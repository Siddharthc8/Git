module top
    
    `include "test_lib.sv"

    initial begin
        run_test("apb_base_test");
    end
    

endmodule 
