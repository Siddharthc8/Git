`timescale 1ns / 1ps




module a30_977_Squares_of_a_Sorted_Array();


endmodule