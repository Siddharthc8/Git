`timescale 1ns / 1ps




module single_port_sync_sram_with_decoder_structural();


endmodule