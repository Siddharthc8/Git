`timescale 1ns / 1ps




module a27_49_Group_Anagrams();


endmodule