`timescale 1ns / 1ps




module a31_344_Reverse_String();


endmodule