`timescale 1ns / 1ps




module a36_16_3Sum_Closest();


endmodule