`timescale 1ns / 1ps




module a33_125_Valid_Palindrome();


endmodule