`timescale 1ns / 1ps




module tb_single_port_sync_sram_behav();


endmodule