`timescale 1ns / 1ps




module a32_167_Two_Sum_II_Input_Array_Is_Sorted();


endmodule