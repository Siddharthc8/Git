`timescale 1ns / 1ps




module tb_detect_pattern_fsm();


endmodule