`timescale 1ns / 1ps




module tb_option_vs_type_option();


endmodule