`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/12/2025 11:21:51 AM
// Design Name: 
// Module Name: tb_kill_task
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_kill_task();


// tasklist | findstr xsim    // To find the tasks list

//  taskkill /F /IM xsimk.exe   // To kill the tasks
endmodule
