input [2:0] a, b,
  input rst,
  input feed,
  output [2:0] y,
  output done

