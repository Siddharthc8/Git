`timescale 1ns/1ps

module tb_assignments();

	tb_a31 a31();
	tb_a32 a32();
	tb_a33 a33();
	tb_a34 a34();
	tb_a35 a35();
	tb_a51 a51();
	tb_a52 a52();
	tb_a53 a53();
	tb_a54 a54();
	tb_a55 a55();
	tb_a56 a56();
	tb_a57 a57();
	tb_a61 a61();
	tb_a62 a62();
	tb_a63 a63();
	tb_a64 a64();
	tb_a65 a65();
	tb_a81 a81();
	
endmodule