`timescale 1ns / 1ps




module reg_file_2_read_1_write_behav();


endmodule