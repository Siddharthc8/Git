`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/10/2024 10:11:29 PM
// Design Name: 
// Module Name: tb_arrays
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_arrays();

    tb_arrays_in_sv a1();
    tb_copying_arrays a2();
    tb_compare_arrays a3();
    tb_dynamic_array a4();
//    tb_a31 e1();
    
endmodule
