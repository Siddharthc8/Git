`timescale 1ns / 1ps




module detect_pattern_fsm();


endmodule